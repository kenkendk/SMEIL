library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

--library SYSTEM_TYPES;
use work.SYSTEM_TYPES.ALL;

--library CUSTOM_TYPES;
use work.CUSTOM_TYPES.ALL;

-- User defined packages here
-- #### USER-DATA-IMPORTS-START
-- #### USER-DATA-IMPORTS-END
entity plusone is
    port(
        -- Bus plusout signals
        plusout_val: out SIGNED(31 DOWNTO 0);
        -- Bus idout signals
        inbus_val: in SIGNED(31 DOWNTO 0);

        -- User defined signals here
        -- #### USER-DATA-ENTITYSIGNALS-START
        -- #### USER-DATA-ENTITYSIGNALS-END

        -- Clock signal
        CLK : in Std_logic;

        --Ready signal
        RDY : in Std_logic;

        --Finished signal
        FIN : out Std_logic;

        --Enable signal
        ENB : in Std_logic;

        --Reset signal
        RST : in Std_logic
    );
end plusone;

architecture RTL of plusone is
    -- User defined signals here
    -- #### USER-DATA-SIGNALS-START
    -- #### USER-DATA-SIGNALS-END

begin

    -- Custom processes go here
    -- #### USER-DATA-PROCESSES-START
    -- #### USER-DATA-PROCESSES-END

    process(

        --Custom sensitivity signals here
        -- #### USER-DATA-SENSITIVITY-START
        -- #### USER-DATA-SENSITIVITY-END

        RDY,
        RST

    )
    variable reentry_guard: std_logic;

    -- #### USER-DATA-NONCLOCKEDVARIABLES-START
    -- #### USER-DATA-NONCLOCKEDVARIABLES-END

    begin
        --Initialize code here
        -- #### USER-DATA-NONCLOCKEDSHAREDINITIALIZECODE-START
        -- #### USER-DATA-NONCLOCKEDSHAREDINITIALIZECODE-END

        if RST = '1' then
            reentry_guard := '0';
            FIN <= '0';

            --Initialize code here
            -- #### USER-DATA-NONCLOCKEDRESETCODE-START
            -- #### USER-DATA-NONCLOCKEDRESETCODE-END

        elsif reentry_guard /= RDY then

            plusout_val <= inbus_val + (1);
            reentry_guard:= RDY;

            --Initialize code here
            -- #### USER-DATA-NONCLOCKEDINITIALIZECODE-START
            -- #### USER-DATA-NONCLOCKEDINITIALIZECODE-END

            FIN <= RDY;
        end if;
    end process;
end RTL;

--User defined architectures here
-- #### USER-DATA-ARCH-START
-- #### USER-DATA-ARCH-END

